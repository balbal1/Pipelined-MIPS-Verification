module pipelined_mips_sva (pipelined_mips_if.DUT _if);
    
endmodule
