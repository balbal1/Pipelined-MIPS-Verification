module pipelined_mips(pipelined_mips_if.DUT _if);
    
    bit [31:0] instruction_memory [0:1023];
    bit [31:0] data_memory [0:1023];

endmodule
